.source quad.net
